---------------------------------------------------------------------------
-- RISC-V-LITE top level entity
---------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity risc_v_dp is
	port
	(	
		
	);